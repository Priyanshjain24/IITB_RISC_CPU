library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Adder is
  port (
    A: in std_logic_vector(15 downto 0);   
    C: out std_logic_vector(15 downto 0)    
  );
end Adder;

architecture Behavioral of Adder is
begin
  C <= std_logic_vector(unsigned(A) + 2);  
end Behavioral;